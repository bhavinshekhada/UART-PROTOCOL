module led(input i_Clock ,input a, output b);
reg b;
parameter clk_cycle9600 = 2500000;
parameter clk_cycle19200 = 5000000;
parameter clk_cycle38400 = 7500000;
parameter clk_cycle57600 = 10000000;
